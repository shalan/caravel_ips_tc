magic
tech sky130A
magscale 1 2
timestamp 1686236622
<< obsli1 >>
rect 1104 2159 120888 491793
<< obsm1 >>
rect 934 1164 120888 491824
<< metal2 >>
rect 2962 0 3018 800
rect 4066 0 4122 800
rect 5170 0 5226 800
rect 6274 0 6330 800
rect 7378 0 7434 800
rect 8482 0 8538 800
rect 9586 0 9642 800
rect 10690 0 10746 800
rect 11794 0 11850 800
rect 12898 0 12954 800
rect 14002 0 14058 800
rect 15106 0 15162 800
rect 16210 0 16266 800
rect 17314 0 17370 800
rect 18418 0 18474 800
rect 19522 0 19578 800
rect 20626 0 20682 800
rect 21730 0 21786 800
rect 22834 0 22890 800
rect 23938 0 23994 800
rect 25042 0 25098 800
rect 26146 0 26202 800
rect 27250 0 27306 800
rect 28354 0 28410 800
rect 29458 0 29514 800
rect 30562 0 30618 800
rect 31666 0 31722 800
rect 32770 0 32826 800
rect 33874 0 33930 800
rect 34978 0 35034 800
rect 36082 0 36138 800
rect 37186 0 37242 800
rect 38290 0 38346 800
rect 39394 0 39450 800
rect 40498 0 40554 800
rect 41602 0 41658 800
rect 42706 0 42762 800
rect 43810 0 43866 800
rect 44914 0 44970 800
rect 46018 0 46074 800
rect 47122 0 47178 800
rect 48226 0 48282 800
rect 49330 0 49386 800
rect 50434 0 50490 800
rect 51538 0 51594 800
rect 52642 0 52698 800
rect 53746 0 53802 800
rect 54850 0 54906 800
rect 55954 0 56010 800
rect 57058 0 57114 800
rect 58162 0 58218 800
rect 59266 0 59322 800
rect 60370 0 60426 800
rect 61474 0 61530 800
rect 62578 0 62634 800
rect 63682 0 63738 800
rect 64786 0 64842 800
rect 65890 0 65946 800
rect 66994 0 67050 800
rect 68098 0 68154 800
rect 69202 0 69258 800
rect 70306 0 70362 800
rect 71410 0 71466 800
rect 72514 0 72570 800
rect 73618 0 73674 800
rect 74722 0 74778 800
rect 75826 0 75882 800
rect 76930 0 76986 800
rect 78034 0 78090 800
rect 79138 0 79194 800
rect 80242 0 80298 800
rect 81346 0 81402 800
rect 82450 0 82506 800
rect 83554 0 83610 800
rect 84658 0 84714 800
rect 85762 0 85818 800
rect 86866 0 86922 800
rect 87970 0 88026 800
rect 89074 0 89130 800
rect 90178 0 90234 800
rect 91282 0 91338 800
rect 92386 0 92442 800
rect 93490 0 93546 800
rect 94594 0 94650 800
rect 95698 0 95754 800
rect 96802 0 96858 800
rect 97906 0 97962 800
rect 99010 0 99066 800
rect 100114 0 100170 800
rect 101218 0 101274 800
rect 102322 0 102378 800
rect 103426 0 103482 800
rect 104530 0 104586 800
rect 105634 0 105690 800
rect 106738 0 106794 800
rect 107842 0 107898 800
rect 108946 0 109002 800
rect 110050 0 110106 800
rect 111154 0 111210 800
rect 112258 0 112314 800
rect 113362 0 113418 800
rect 114466 0 114522 800
rect 115570 0 115626 800
rect 116674 0 116730 800
rect 117778 0 117834 800
rect 118882 0 118938 800
<< obsm2 >>
rect 938 856 120594 491813
rect 938 734 2906 856
rect 3074 734 4010 856
rect 4178 734 5114 856
rect 5282 734 6218 856
rect 6386 734 7322 856
rect 7490 734 8426 856
rect 8594 734 9530 856
rect 9698 734 10634 856
rect 10802 734 11738 856
rect 11906 734 12842 856
rect 13010 734 13946 856
rect 14114 734 15050 856
rect 15218 734 16154 856
rect 16322 734 17258 856
rect 17426 734 18362 856
rect 18530 734 19466 856
rect 19634 734 20570 856
rect 20738 734 21674 856
rect 21842 734 22778 856
rect 22946 734 23882 856
rect 24050 734 24986 856
rect 25154 734 26090 856
rect 26258 734 27194 856
rect 27362 734 28298 856
rect 28466 734 29402 856
rect 29570 734 30506 856
rect 30674 734 31610 856
rect 31778 734 32714 856
rect 32882 734 33818 856
rect 33986 734 34922 856
rect 35090 734 36026 856
rect 36194 734 37130 856
rect 37298 734 38234 856
rect 38402 734 39338 856
rect 39506 734 40442 856
rect 40610 734 41546 856
rect 41714 734 42650 856
rect 42818 734 43754 856
rect 43922 734 44858 856
rect 45026 734 45962 856
rect 46130 734 47066 856
rect 47234 734 48170 856
rect 48338 734 49274 856
rect 49442 734 50378 856
rect 50546 734 51482 856
rect 51650 734 52586 856
rect 52754 734 53690 856
rect 53858 734 54794 856
rect 54962 734 55898 856
rect 56066 734 57002 856
rect 57170 734 58106 856
rect 58274 734 59210 856
rect 59378 734 60314 856
rect 60482 734 61418 856
rect 61586 734 62522 856
rect 62690 734 63626 856
rect 63794 734 64730 856
rect 64898 734 65834 856
rect 66002 734 66938 856
rect 67106 734 68042 856
rect 68210 734 69146 856
rect 69314 734 70250 856
rect 70418 734 71354 856
rect 71522 734 72458 856
rect 72626 734 73562 856
rect 73730 734 74666 856
rect 74834 734 75770 856
rect 75938 734 76874 856
rect 77042 734 77978 856
rect 78146 734 79082 856
rect 79250 734 80186 856
rect 80354 734 81290 856
rect 81458 734 82394 856
rect 82562 734 83498 856
rect 83666 734 84602 856
rect 84770 734 85706 856
rect 85874 734 86810 856
rect 86978 734 87914 856
rect 88082 734 89018 856
rect 89186 734 90122 856
rect 90290 734 91226 856
rect 91394 734 92330 856
rect 92498 734 93434 856
rect 93602 734 94538 856
rect 94706 734 95642 856
rect 95810 734 96746 856
rect 96914 734 97850 856
rect 98018 734 98954 856
rect 99122 734 100058 856
rect 100226 734 101162 856
rect 101330 734 102266 856
rect 102434 734 103370 856
rect 103538 734 104474 856
rect 104642 734 105578 856
rect 105746 734 106682 856
rect 106850 734 107786 856
rect 107954 734 108890 856
rect 109058 734 109994 856
rect 110162 734 111098 856
rect 111266 734 112202 856
rect 112370 734 113306 856
rect 113474 734 114410 856
rect 114578 734 115514 856
rect 115682 734 116618 856
rect 116786 734 117722 856
rect 117890 734 118826 856
rect 118994 734 120594 856
<< metal3 >>
rect 0 483352 800 483472
rect 0 467032 800 467152
rect 0 450712 800 450832
rect 0 434392 800 434512
rect 0 418072 800 418192
rect 0 401752 800 401872
rect 0 385432 800 385552
rect 0 369112 800 369232
rect 0 352792 800 352912
rect 0 336472 800 336592
rect 0 320152 800 320272
rect 0 303832 800 303952
rect 0 287512 800 287632
rect 0 271192 800 271312
rect 0 254872 800 254992
rect 0 238552 800 238672
rect 0 222232 800 222352
rect 0 205912 800 206032
rect 0 189592 800 189712
rect 0 173272 800 173392
rect 0 156952 800 157072
rect 0 140632 800 140752
rect 0 124312 800 124432
rect 0 107992 800 108112
rect 0 91672 800 91792
rect 0 75352 800 75472
rect 0 59032 800 59152
rect 0 42712 800 42832
rect 0 26392 800 26512
rect 121200 24760 122000 24880
rect 121200 15512 122000 15632
rect 0 10072 800 10192
rect 121200 6264 122000 6384
<< obsm3 >>
rect 800 483552 121200 491809
rect 880 483272 121200 483552
rect 800 467232 121200 483272
rect 880 466952 121200 467232
rect 800 450912 121200 466952
rect 880 450632 121200 450912
rect 800 434592 121200 450632
rect 880 434312 121200 434592
rect 800 418272 121200 434312
rect 880 417992 121200 418272
rect 800 401952 121200 417992
rect 880 401672 121200 401952
rect 800 385632 121200 401672
rect 880 385352 121200 385632
rect 800 369312 121200 385352
rect 880 369032 121200 369312
rect 800 352992 121200 369032
rect 880 352712 121200 352992
rect 800 336672 121200 352712
rect 880 336392 121200 336672
rect 800 320352 121200 336392
rect 880 320072 121200 320352
rect 800 304032 121200 320072
rect 880 303752 121200 304032
rect 800 287712 121200 303752
rect 880 287432 121200 287712
rect 800 271392 121200 287432
rect 880 271112 121200 271392
rect 800 255072 121200 271112
rect 880 254792 121200 255072
rect 800 238752 121200 254792
rect 880 238472 121200 238752
rect 800 222432 121200 238472
rect 880 222152 121200 222432
rect 800 206112 121200 222152
rect 880 205832 121200 206112
rect 800 189792 121200 205832
rect 880 189512 121200 189792
rect 800 173472 121200 189512
rect 880 173192 121200 173472
rect 800 157152 121200 173192
rect 880 156872 121200 157152
rect 800 140832 121200 156872
rect 880 140552 121200 140832
rect 800 124512 121200 140552
rect 880 124232 121200 124512
rect 800 108192 121200 124232
rect 880 107912 121200 108192
rect 800 91872 121200 107912
rect 880 91592 121200 91872
rect 800 75552 121200 91592
rect 880 75272 121200 75552
rect 800 59232 121200 75272
rect 880 58952 121200 59232
rect 800 42912 121200 58952
rect 880 42632 121200 42912
rect 800 26592 121200 42632
rect 880 26312 121200 26592
rect 800 24960 121200 26312
rect 800 24680 121120 24960
rect 800 15712 121200 24680
rect 800 15432 121120 15712
rect 800 10272 121200 15432
rect 880 9992 121200 10272
rect 800 6464 121200 9992
rect 800 6184 121120 6464
rect 800 1803 121200 6184
<< metal4 >>
rect 4048 2128 4688 491824
rect 12208 2128 12848 491824
rect 20368 2128 21008 491824
rect 28528 2128 29168 491824
rect 36688 2128 37328 491824
rect 44848 2128 45488 491824
rect 53008 2128 53648 491824
rect 61168 2128 61808 491824
rect 69328 2128 69968 491824
rect 77488 2128 78128 491824
rect 85648 2128 86288 491824
rect 93808 2128 94448 491824
rect 101968 2128 102608 491824
rect 110128 2128 110768 491824
rect 118288 2128 118928 491824
<< obsm4 >>
rect 22507 2347 28448 161941
rect 29248 2347 36608 161941
rect 37408 2347 44768 161941
rect 45568 2347 52928 161941
rect 53728 2347 61088 161941
rect 61888 2347 69248 161941
rect 70048 2347 77408 161941
rect 78208 2347 84397 161941
<< labels >>
rlabel metal4 s 110128 2128 110768 491824 6 VGND
port 1 nsew ground default
rlabel metal4 s 93808 2128 94448 491824 6 VGND
port 1 nsew ground default
rlabel metal4 s 77488 2128 78128 491824 6 VGND
port 1 nsew ground default
rlabel metal4 s 61168 2128 61808 491824 6 VGND
port 1 nsew ground default
rlabel metal4 s 44848 2128 45488 491824 6 VGND
port 1 nsew ground default
rlabel metal4 s 28528 2128 29168 491824 6 VGND
port 1 nsew ground default
rlabel metal4 s 12208 2128 12848 491824 6 VGND
port 1 nsew ground default
rlabel metal4 s 118288 2128 118928 491824 6 VPWR
port 2 nsew power default
rlabel metal4 s 101968 2128 102608 491824 6 VPWR
port 2 nsew power default
rlabel metal4 s 85648 2128 86288 491824 6 VPWR
port 2 nsew power default
rlabel metal4 s 69328 2128 69968 491824 6 VPWR
port 2 nsew power default
rlabel metal4 s 53008 2128 53648 491824 6 VPWR
port 2 nsew power default
rlabel metal4 s 36688 2128 37328 491824 6 VPWR
port 2 nsew power default
rlabel metal4 s 20368 2128 21008 491824 6 VPWR
port 2 nsew power default
rlabel metal4 s 4048 2128 4688 491824 6 VPWR
port 2 nsew power default
rlabel metal3 s 0 483352 800 483472 6 io_in[0]
port 3 nsew
rlabel metal3 s 0 434392 800 434512 6 io_in[1]
port 4 nsew
rlabel metal3 s 0 385432 800 385552 6 io_in[2]
port 5 nsew
rlabel metal3 s 0 336472 800 336592 6 io_in[3]
port 6 nsew
rlabel metal3 s 0 287512 800 287632 6 io_in[4]
port 7 nsew
rlabel metal3 s 0 238552 800 238672 6 io_in[5]
port 8 nsew
rlabel metal3 s 0 189592 800 189712 6 io_in[6]
port 9 nsew
rlabel metal3 s 0 140632 800 140752 6 io_in[7]
port 10 nsew
rlabel metal3 s 0 91672 800 91792 6 io_in[8]
port 11 nsew
rlabel metal3 s 0 42712 800 42832 6 io_in[9]
port 12 nsew
rlabel metal3 s 0 450712 800 450832 6 io_oeb[0]
port 13 nsew
rlabel metal3 s 0 401752 800 401872 6 io_oeb[1]
port 14 nsew
rlabel metal3 s 0 352792 800 352912 6 io_oeb[2]
port 15 nsew
rlabel metal3 s 0 303832 800 303952 6 io_oeb[3]
port 16 nsew
rlabel metal3 s 0 254872 800 254992 6 io_oeb[4]
port 17 nsew
rlabel metal3 s 0 205912 800 206032 6 io_oeb[5]
port 18 nsew
rlabel metal3 s 0 156952 800 157072 6 io_oeb[6]
port 19 nsew
rlabel metal3 s 0 107992 800 108112 6 io_oeb[7]
port 20 nsew
rlabel metal3 s 0 59032 800 59152 6 io_oeb[8]
port 21 nsew
rlabel metal3 s 0 10072 800 10192 6 io_oeb[9]
port 22 nsew
rlabel metal3 s 0 467032 800 467152 6 io_out[0]
port 23 nsew
rlabel metal3 s 0 418072 800 418192 6 io_out[1]
port 24 nsew
rlabel metal3 s 0 369112 800 369232 6 io_out[2]
port 25 nsew
rlabel metal3 s 0 320152 800 320272 6 io_out[3]
port 26 nsew
rlabel metal3 s 0 271192 800 271312 6 io_out[4]
port 27 nsew
rlabel metal3 s 0 222232 800 222352 6 io_out[5]
port 28 nsew
rlabel metal3 s 0 173272 800 173392 6 io_out[6]
port 29 nsew
rlabel metal3 s 0 124312 800 124432 6 io_out[7]
port 30 nsew
rlabel metal3 s 0 75352 800 75472 6 io_out[8]
port 31 nsew
rlabel metal3 s 0 26392 800 26512 6 io_out[9]
port 32 nsew
rlabel metal3 s 121200 6264 122000 6384 6 irq[0]
port 33 nsew
rlabel metal3 s 121200 15512 122000 15632 6 irq[1]
port 34 nsew
rlabel metal3 s 121200 24760 122000 24880 6 irq[2]
port 35 nsew
rlabel metal2 s 2962 0 3018 800 6 wb_clk_i
port 36 nsew
rlabel metal2 s 4066 0 4122 800 6 wb_rst_i
port 37 nsew
rlabel metal2 s 5170 0 5226 800 6 wbs_ack_o
port 38 nsew
rlabel metal2 s 9586 0 9642 800 6 wbs_adr_i[0]
port 39 nsew
rlabel metal2 s 47122 0 47178 800 6 wbs_adr_i[10]
port 40 nsew
rlabel metal2 s 50434 0 50490 800 6 wbs_adr_i[11]
port 41 nsew
rlabel metal2 s 53746 0 53802 800 6 wbs_adr_i[12]
port 42 nsew
rlabel metal2 s 57058 0 57114 800 6 wbs_adr_i[13]
port 43 nsew
rlabel metal2 s 60370 0 60426 800 6 wbs_adr_i[14]
port 44 nsew
rlabel metal2 s 63682 0 63738 800 6 wbs_adr_i[15]
port 45 nsew
rlabel metal2 s 66994 0 67050 800 6 wbs_adr_i[16]
port 46 nsew
rlabel metal2 s 70306 0 70362 800 6 wbs_adr_i[17]
port 47 nsew
rlabel metal2 s 73618 0 73674 800 6 wbs_adr_i[18]
port 48 nsew
rlabel metal2 s 76930 0 76986 800 6 wbs_adr_i[19]
port 49 nsew
rlabel metal2 s 14002 0 14058 800 6 wbs_adr_i[1]
port 50 nsew
rlabel metal2 s 80242 0 80298 800 6 wbs_adr_i[20]
port 51 nsew
rlabel metal2 s 83554 0 83610 800 6 wbs_adr_i[21]
port 52 nsew
rlabel metal2 s 86866 0 86922 800 6 wbs_adr_i[22]
port 53 nsew
rlabel metal2 s 90178 0 90234 800 6 wbs_adr_i[23]
port 54 nsew
rlabel metal2 s 93490 0 93546 800 6 wbs_adr_i[24]
port 55 nsew
rlabel metal2 s 96802 0 96858 800 6 wbs_adr_i[25]
port 56 nsew
rlabel metal2 s 100114 0 100170 800 6 wbs_adr_i[26]
port 57 nsew
rlabel metal2 s 103426 0 103482 800 6 wbs_adr_i[27]
port 58 nsew
rlabel metal2 s 106738 0 106794 800 6 wbs_adr_i[28]
port 59 nsew
rlabel metal2 s 110050 0 110106 800 6 wbs_adr_i[29]
port 60 nsew
rlabel metal2 s 18418 0 18474 800 6 wbs_adr_i[2]
port 61 nsew
rlabel metal2 s 113362 0 113418 800 6 wbs_adr_i[30]
port 62 nsew
rlabel metal2 s 116674 0 116730 800 6 wbs_adr_i[31]
port 63 nsew
rlabel metal2 s 22834 0 22890 800 6 wbs_adr_i[3]
port 64 nsew
rlabel metal2 s 27250 0 27306 800 6 wbs_adr_i[4]
port 65 nsew
rlabel metal2 s 30562 0 30618 800 6 wbs_adr_i[5]
port 66 nsew
rlabel metal2 s 33874 0 33930 800 6 wbs_adr_i[6]
port 67 nsew
rlabel metal2 s 37186 0 37242 800 6 wbs_adr_i[7]
port 68 nsew
rlabel metal2 s 40498 0 40554 800 6 wbs_adr_i[8]
port 69 nsew
rlabel metal2 s 43810 0 43866 800 6 wbs_adr_i[9]
port 70 nsew
rlabel metal2 s 6274 0 6330 800 6 wbs_cyc_i
port 71 nsew
rlabel metal2 s 10690 0 10746 800 6 wbs_dat_i[0]
port 72 nsew
rlabel metal2 s 48226 0 48282 800 6 wbs_dat_i[10]
port 73 nsew
rlabel metal2 s 51538 0 51594 800 6 wbs_dat_i[11]
port 74 nsew
rlabel metal2 s 54850 0 54906 800 6 wbs_dat_i[12]
port 75 nsew
rlabel metal2 s 58162 0 58218 800 6 wbs_dat_i[13]
port 76 nsew
rlabel metal2 s 61474 0 61530 800 6 wbs_dat_i[14]
port 77 nsew
rlabel metal2 s 64786 0 64842 800 6 wbs_dat_i[15]
port 78 nsew
rlabel metal2 s 68098 0 68154 800 6 wbs_dat_i[16]
port 79 nsew
rlabel metal2 s 71410 0 71466 800 6 wbs_dat_i[17]
port 80 nsew
rlabel metal2 s 74722 0 74778 800 6 wbs_dat_i[18]
port 81 nsew
rlabel metal2 s 78034 0 78090 800 6 wbs_dat_i[19]
port 82 nsew
rlabel metal2 s 15106 0 15162 800 6 wbs_dat_i[1]
port 83 nsew
rlabel metal2 s 81346 0 81402 800 6 wbs_dat_i[20]
port 84 nsew
rlabel metal2 s 84658 0 84714 800 6 wbs_dat_i[21]
port 85 nsew
rlabel metal2 s 87970 0 88026 800 6 wbs_dat_i[22]
port 86 nsew
rlabel metal2 s 91282 0 91338 800 6 wbs_dat_i[23]
port 87 nsew
rlabel metal2 s 94594 0 94650 800 6 wbs_dat_i[24]
port 88 nsew
rlabel metal2 s 97906 0 97962 800 6 wbs_dat_i[25]
port 89 nsew
rlabel metal2 s 101218 0 101274 800 6 wbs_dat_i[26]
port 90 nsew
rlabel metal2 s 104530 0 104586 800 6 wbs_dat_i[27]
port 91 nsew
rlabel metal2 s 107842 0 107898 800 6 wbs_dat_i[28]
port 92 nsew
rlabel metal2 s 111154 0 111210 800 6 wbs_dat_i[29]
port 93 nsew
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_i[2]
port 94 nsew
rlabel metal2 s 114466 0 114522 800 6 wbs_dat_i[30]
port 95 nsew
rlabel metal2 s 117778 0 117834 800 6 wbs_dat_i[31]
port 96 nsew
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_i[3]
port 97 nsew
rlabel metal2 s 28354 0 28410 800 6 wbs_dat_i[4]
port 98 nsew
rlabel metal2 s 31666 0 31722 800 6 wbs_dat_i[5]
port 99 nsew
rlabel metal2 s 34978 0 35034 800 6 wbs_dat_i[6]
port 100 nsew
rlabel metal2 s 38290 0 38346 800 6 wbs_dat_i[7]
port 101 nsew
rlabel metal2 s 41602 0 41658 800 6 wbs_dat_i[8]
port 102 nsew
rlabel metal2 s 44914 0 44970 800 6 wbs_dat_i[9]
port 103 nsew
rlabel metal2 s 11794 0 11850 800 6 wbs_dat_o[0]
port 104 nsew
rlabel metal2 s 49330 0 49386 800 6 wbs_dat_o[10]
port 105 nsew
rlabel metal2 s 52642 0 52698 800 6 wbs_dat_o[11]
port 106 nsew
rlabel metal2 s 55954 0 56010 800 6 wbs_dat_o[12]
port 107 nsew
rlabel metal2 s 59266 0 59322 800 6 wbs_dat_o[13]
port 108 nsew
rlabel metal2 s 62578 0 62634 800 6 wbs_dat_o[14]
port 109 nsew
rlabel metal2 s 65890 0 65946 800 6 wbs_dat_o[15]
port 110 nsew
rlabel metal2 s 69202 0 69258 800 6 wbs_dat_o[16]
port 111 nsew
rlabel metal2 s 72514 0 72570 800 6 wbs_dat_o[17]
port 112 nsew
rlabel metal2 s 75826 0 75882 800 6 wbs_dat_o[18]
port 113 nsew
rlabel metal2 s 79138 0 79194 800 6 wbs_dat_o[19]
port 114 nsew
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_o[1]
port 115 nsew
rlabel metal2 s 82450 0 82506 800 6 wbs_dat_o[20]
port 116 nsew
rlabel metal2 s 85762 0 85818 800 6 wbs_dat_o[21]
port 117 nsew
rlabel metal2 s 89074 0 89130 800 6 wbs_dat_o[22]
port 118 nsew
rlabel metal2 s 92386 0 92442 800 6 wbs_dat_o[23]
port 119 nsew
rlabel metal2 s 95698 0 95754 800 6 wbs_dat_o[24]
port 120 nsew
rlabel metal2 s 99010 0 99066 800 6 wbs_dat_o[25]
port 121 nsew
rlabel metal2 s 102322 0 102378 800 6 wbs_dat_o[26]
port 122 nsew
rlabel metal2 s 105634 0 105690 800 6 wbs_dat_o[27]
port 123 nsew
rlabel metal2 s 108946 0 109002 800 6 wbs_dat_o[28]
port 124 nsew
rlabel metal2 s 112258 0 112314 800 6 wbs_dat_o[29]
port 125 nsew
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_o[2]
port 126 nsew
rlabel metal2 s 115570 0 115626 800 6 wbs_dat_o[30]
port 127 nsew
rlabel metal2 s 118882 0 118938 800 6 wbs_dat_o[31]
port 128 nsew
rlabel metal2 s 25042 0 25098 800 6 wbs_dat_o[3]
port 129 nsew
rlabel metal2 s 29458 0 29514 800 6 wbs_dat_o[4]
port 130 nsew
rlabel metal2 s 32770 0 32826 800 6 wbs_dat_o[5]
port 131 nsew
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_o[6]
port 132 nsew
rlabel metal2 s 39394 0 39450 800 6 wbs_dat_o[7]
port 133 nsew
rlabel metal2 s 42706 0 42762 800 6 wbs_dat_o[8]
port 134 nsew
rlabel metal2 s 46018 0 46074 800 6 wbs_dat_o[9]
port 135 nsew
rlabel metal2 s 12898 0 12954 800 6 wbs_sel_i[0]
port 136 nsew
rlabel metal2 s 17314 0 17370 800 6 wbs_sel_i[1]
port 137 nsew
rlabel metal2 s 21730 0 21786 800 6 wbs_sel_i[2]
port 138 nsew
rlabel metal2 s 26146 0 26202 800 6 wbs_sel_i[3]
port 139 nsew
rlabel metal2 s 7378 0 7434 800 6 wbs_stb_i
port 140 nsew
rlabel metal2 s 8482 0 8538 800 6 wbs_we_i
port 141 nsew
<< properties >>
string FIXED_BBOX 0 0 122000 494000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 38579772
string GDS_FILE /home/hosni/caravel_ips/caravel_ips_tc/openlane/caravel_ips/runs/23_06_08_07_55/results/signoff/caravel_ips.magic.gds
string GDS_START 1121362
<< end >>

