VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravel_ips
  CLASS BLOCK ;
  FOREIGN caravel_ips ;
  ORIGIN 0.000 0.000 ;
  SIZE 610.000 BY 2470.000 ;
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 550.640 10.640 553.840 2459.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 469.040 10.640 472.240 2459.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.440 10.640 390.640 2459.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 305.840 10.640 309.040 2459.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 224.240 10.640 227.440 2459.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 142.640 10.640 145.840 2459.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 61.040 10.640 64.240 2459.120 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 591.440 10.640 594.640 2459.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 509.840 10.640 513.040 2459.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 428.240 10.640 431.440 2459.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.640 10.640 349.840 2459.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 265.040 10.640 268.240 2459.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 183.440 10.640 186.640 2459.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 101.840 10.640 105.040 2459.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 20.240 10.640 23.440 2459.120 ;
    END
  END VPWR
  PIN io_in[0]
    PORT
      LAYER met3 ;
        RECT 0.000 2416.760 4.000 2417.360 ;
    END
  END io_in[0]
  PIN io_in[1]
    PORT
      LAYER met3 ;
        RECT 0.000 2171.960 4.000 2172.560 ;
    END
  END io_in[1]
  PIN io_in[2]
    PORT
      LAYER met3 ;
        RECT 0.000 1927.160 4.000 1927.760 ;
    END
  END io_in[2]
  PIN io_in[3]
    PORT
      LAYER met3 ;
        RECT 0.000 1682.360 4.000 1682.960 ;
    END
  END io_in[3]
  PIN io_in[4]
    PORT
      LAYER met3 ;
        RECT 0.000 1437.560 4.000 1438.160 ;
    END
  END io_in[4]
  PIN io_in[5]
    PORT
      LAYER met3 ;
        RECT 0.000 1192.760 4.000 1193.360 ;
    END
  END io_in[5]
  PIN io_in[6]
    PORT
      LAYER met3 ;
        RECT 0.000 947.960 4.000 948.560 ;
    END
  END io_in[6]
  PIN io_in[7]
    PORT
      LAYER met3 ;
        RECT 0.000 703.160 4.000 703.760 ;
    END
  END io_in[7]
  PIN io_in[8]
    PORT
      LAYER met3 ;
        RECT 0.000 458.360 4.000 458.960 ;
    END
  END io_in[8]
  PIN io_in[9]
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    PORT
      LAYER met3 ;
        RECT 0.000 2253.560 4.000 2254.160 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    PORT
      LAYER met3 ;
        RECT 0.000 2008.760 4.000 2009.360 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    PORT
      LAYER met3 ;
        RECT 0.000 1763.960 4.000 1764.560 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    PORT
      LAYER met3 ;
        RECT 0.000 1519.160 4.000 1519.760 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    PORT
      LAYER met3 ;
        RECT 0.000 1274.360 4.000 1274.960 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    PORT
      LAYER met3 ;
        RECT 0.000 1029.560 4.000 1030.160 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    PORT
      LAYER met3 ;
        RECT 0.000 784.760 4.000 785.360 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    PORT
      LAYER met3 ;
        RECT 0.000 539.960 4.000 540.560 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    PORT
      LAYER met3 ;
        RECT 0.000 2335.160 4.000 2335.760 ;
    END
  END io_out[0]
  PIN io_out[1]
    PORT
      LAYER met3 ;
        RECT 0.000 2090.360 4.000 2090.960 ;
    END
  END io_out[1]
  PIN io_out[2]
    PORT
      LAYER met3 ;
        RECT 0.000 1845.560 4.000 1846.160 ;
    END
  END io_out[2]
  PIN io_out[3]
    PORT
      LAYER met3 ;
        RECT 0.000 1600.760 4.000 1601.360 ;
    END
  END io_out[3]
  PIN io_out[4]
    PORT
      LAYER met3 ;
        RECT 0.000 1355.960 4.000 1356.560 ;
    END
  END io_out[4]
  PIN io_out[5]
    PORT
      LAYER met3 ;
        RECT 0.000 1111.160 4.000 1111.760 ;
    END
  END io_out[5]
  PIN io_out[6]
    PORT
      LAYER met3 ;
        RECT 0.000 866.360 4.000 866.960 ;
    END
  END io_out[6]
  PIN io_out[7]
    PORT
      LAYER met3 ;
        RECT 0.000 621.560 4.000 622.160 ;
    END
  END io_out[7]
  PIN io_out[8]
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END io_out[8]
  PIN io_out[9]
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END io_out[9]
  PIN irq[0]
    PORT
      LAYER met3 ;
        RECT 606.000 31.320 610.000 31.920 ;
    END
  END irq[0]
  PIN irq[1]
    PORT
      LAYER met3 ;
        RECT 606.000 77.560 610.000 78.160 ;
    END
  END irq[1]
  PIN irq[2]
    PORT
      LAYER met3 ;
        RECT 606.000 123.800 610.000 124.400 ;
    END
  END irq[2]
  PIN wb_clk_i
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    PORT
      LAYER met2 ;
        RECT 268.730 0.000 269.010 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    PORT
      LAYER met2 ;
        RECT 351.530 0.000 351.810 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    PORT
      LAYER met2 ;
        RECT 384.650 0.000 384.930 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    PORT
      LAYER met2 ;
        RECT 401.210 0.000 401.490 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    PORT
      LAYER met2 ;
        RECT 417.770 0.000 418.050 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    PORT
      LAYER met2 ;
        RECT 434.330 0.000 434.610 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    PORT
      LAYER met2 ;
        RECT 467.450 0.000 467.730 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    PORT
      LAYER met2 ;
        RECT 484.010 0.000 484.290 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    PORT
      LAYER met2 ;
        RECT 500.570 0.000 500.850 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    PORT
      LAYER met2 ;
        RECT 517.130 0.000 517.410 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    PORT
      LAYER met2 ;
        RECT 533.690 0.000 533.970 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    PORT
      LAYER met2 ;
        RECT 550.250 0.000 550.530 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    PORT
      LAYER met2 ;
        RECT 583.370 0.000 583.650 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    PORT
      LAYER met2 ;
        RECT 241.130 0.000 241.410 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    PORT
      LAYER met2 ;
        RECT 290.810 0.000 291.090 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    PORT
      LAYER met2 ;
        RECT 307.370 0.000 307.650 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    PORT
      LAYER met2 ;
        RECT 340.490 0.000 340.770 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    PORT
      LAYER met2 ;
        RECT 390.170 0.000 390.450 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    PORT
      LAYER met2 ;
        RECT 406.730 0.000 407.010 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    PORT
      LAYER met2 ;
        RECT 423.290 0.000 423.570 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    PORT
      LAYER met2 ;
        RECT 439.850 0.000 440.130 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    PORT
      LAYER met2 ;
        RECT 456.410 0.000 456.690 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    PORT
      LAYER met2 ;
        RECT 472.970 0.000 473.250 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    PORT
      LAYER met2 ;
        RECT 506.090 0.000 506.370 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    PORT
      LAYER met2 ;
        RECT 522.650 0.000 522.930 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    PORT
      LAYER met2 ;
        RECT 539.210 0.000 539.490 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    PORT
      LAYER met2 ;
        RECT 555.770 0.000 556.050 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    PORT
      LAYER met2 ;
        RECT 572.330 0.000 572.610 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    PORT
      LAYER met2 ;
        RECT 588.890 0.000 589.170 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    PORT
      LAYER met2 ;
        RECT 263.210 0.000 263.490 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    PORT
      LAYER met2 ;
        RECT 346.010 0.000 346.290 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    PORT
      LAYER met2 ;
        RECT 362.570 0.000 362.850 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    PORT
      LAYER met2 ;
        RECT 428.810 0.000 429.090 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    PORT
      LAYER met2 ;
        RECT 445.370 0.000 445.650 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    PORT
      LAYER met2 ;
        RECT 461.930 0.000 462.210 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    PORT
      LAYER met2 ;
        RECT 478.490 0.000 478.770 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    PORT
      LAYER met2 ;
        RECT 495.050 0.000 495.330 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    PORT
      LAYER met2 ;
        RECT 511.610 0.000 511.890 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    PORT
      LAYER met2 ;
        RECT 544.730 0.000 545.010 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    PORT
      LAYER met2 ;
        RECT 561.290 0.000 561.570 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    PORT
      LAYER met2 ;
        RECT 577.850 0.000 578.130 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    PORT
      LAYER met2 ;
        RECT 594.410 0.000 594.690 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    PORT
      LAYER met2 ;
        RECT 213.530 0.000 213.810 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 604.440 2458.965 ;
      LAYER met1 ;
        RECT 4.670 5.820 604.440 2459.120 ;
      LAYER met2 ;
        RECT 4.690 4.280 602.970 2459.065 ;
        RECT 4.690 3.670 14.530 4.280 ;
        RECT 15.370 3.670 20.050 4.280 ;
        RECT 20.890 3.670 25.570 4.280 ;
        RECT 26.410 3.670 31.090 4.280 ;
        RECT 31.930 3.670 36.610 4.280 ;
        RECT 37.450 3.670 42.130 4.280 ;
        RECT 42.970 3.670 47.650 4.280 ;
        RECT 48.490 3.670 53.170 4.280 ;
        RECT 54.010 3.670 58.690 4.280 ;
        RECT 59.530 3.670 64.210 4.280 ;
        RECT 65.050 3.670 69.730 4.280 ;
        RECT 70.570 3.670 75.250 4.280 ;
        RECT 76.090 3.670 80.770 4.280 ;
        RECT 81.610 3.670 86.290 4.280 ;
        RECT 87.130 3.670 91.810 4.280 ;
        RECT 92.650 3.670 97.330 4.280 ;
        RECT 98.170 3.670 102.850 4.280 ;
        RECT 103.690 3.670 108.370 4.280 ;
        RECT 109.210 3.670 113.890 4.280 ;
        RECT 114.730 3.670 119.410 4.280 ;
        RECT 120.250 3.670 124.930 4.280 ;
        RECT 125.770 3.670 130.450 4.280 ;
        RECT 131.290 3.670 135.970 4.280 ;
        RECT 136.810 3.670 141.490 4.280 ;
        RECT 142.330 3.670 147.010 4.280 ;
        RECT 147.850 3.670 152.530 4.280 ;
        RECT 153.370 3.670 158.050 4.280 ;
        RECT 158.890 3.670 163.570 4.280 ;
        RECT 164.410 3.670 169.090 4.280 ;
        RECT 169.930 3.670 174.610 4.280 ;
        RECT 175.450 3.670 180.130 4.280 ;
        RECT 180.970 3.670 185.650 4.280 ;
        RECT 186.490 3.670 191.170 4.280 ;
        RECT 192.010 3.670 196.690 4.280 ;
        RECT 197.530 3.670 202.210 4.280 ;
        RECT 203.050 3.670 207.730 4.280 ;
        RECT 208.570 3.670 213.250 4.280 ;
        RECT 214.090 3.670 218.770 4.280 ;
        RECT 219.610 3.670 224.290 4.280 ;
        RECT 225.130 3.670 229.810 4.280 ;
        RECT 230.650 3.670 235.330 4.280 ;
        RECT 236.170 3.670 240.850 4.280 ;
        RECT 241.690 3.670 246.370 4.280 ;
        RECT 247.210 3.670 251.890 4.280 ;
        RECT 252.730 3.670 257.410 4.280 ;
        RECT 258.250 3.670 262.930 4.280 ;
        RECT 263.770 3.670 268.450 4.280 ;
        RECT 269.290 3.670 273.970 4.280 ;
        RECT 274.810 3.670 279.490 4.280 ;
        RECT 280.330 3.670 285.010 4.280 ;
        RECT 285.850 3.670 290.530 4.280 ;
        RECT 291.370 3.670 296.050 4.280 ;
        RECT 296.890 3.670 301.570 4.280 ;
        RECT 302.410 3.670 307.090 4.280 ;
        RECT 307.930 3.670 312.610 4.280 ;
        RECT 313.450 3.670 318.130 4.280 ;
        RECT 318.970 3.670 323.650 4.280 ;
        RECT 324.490 3.670 329.170 4.280 ;
        RECT 330.010 3.670 334.690 4.280 ;
        RECT 335.530 3.670 340.210 4.280 ;
        RECT 341.050 3.670 345.730 4.280 ;
        RECT 346.570 3.670 351.250 4.280 ;
        RECT 352.090 3.670 356.770 4.280 ;
        RECT 357.610 3.670 362.290 4.280 ;
        RECT 363.130 3.670 367.810 4.280 ;
        RECT 368.650 3.670 373.330 4.280 ;
        RECT 374.170 3.670 378.850 4.280 ;
        RECT 379.690 3.670 384.370 4.280 ;
        RECT 385.210 3.670 389.890 4.280 ;
        RECT 390.730 3.670 395.410 4.280 ;
        RECT 396.250 3.670 400.930 4.280 ;
        RECT 401.770 3.670 406.450 4.280 ;
        RECT 407.290 3.670 411.970 4.280 ;
        RECT 412.810 3.670 417.490 4.280 ;
        RECT 418.330 3.670 423.010 4.280 ;
        RECT 423.850 3.670 428.530 4.280 ;
        RECT 429.370 3.670 434.050 4.280 ;
        RECT 434.890 3.670 439.570 4.280 ;
        RECT 440.410 3.670 445.090 4.280 ;
        RECT 445.930 3.670 450.610 4.280 ;
        RECT 451.450 3.670 456.130 4.280 ;
        RECT 456.970 3.670 461.650 4.280 ;
        RECT 462.490 3.670 467.170 4.280 ;
        RECT 468.010 3.670 472.690 4.280 ;
        RECT 473.530 3.670 478.210 4.280 ;
        RECT 479.050 3.670 483.730 4.280 ;
        RECT 484.570 3.670 489.250 4.280 ;
        RECT 490.090 3.670 494.770 4.280 ;
        RECT 495.610 3.670 500.290 4.280 ;
        RECT 501.130 3.670 505.810 4.280 ;
        RECT 506.650 3.670 511.330 4.280 ;
        RECT 512.170 3.670 516.850 4.280 ;
        RECT 517.690 3.670 522.370 4.280 ;
        RECT 523.210 3.670 527.890 4.280 ;
        RECT 528.730 3.670 533.410 4.280 ;
        RECT 534.250 3.670 538.930 4.280 ;
        RECT 539.770 3.670 544.450 4.280 ;
        RECT 545.290 3.670 549.970 4.280 ;
        RECT 550.810 3.670 555.490 4.280 ;
        RECT 556.330 3.670 561.010 4.280 ;
        RECT 561.850 3.670 566.530 4.280 ;
        RECT 567.370 3.670 572.050 4.280 ;
        RECT 572.890 3.670 577.570 4.280 ;
        RECT 578.410 3.670 583.090 4.280 ;
        RECT 583.930 3.670 588.610 4.280 ;
        RECT 589.450 3.670 594.130 4.280 ;
        RECT 594.970 3.670 602.970 4.280 ;
      LAYER met3 ;
        RECT 4.000 2417.760 606.000 2459.045 ;
        RECT 4.400 2416.360 606.000 2417.760 ;
        RECT 4.000 2336.160 606.000 2416.360 ;
        RECT 4.400 2334.760 606.000 2336.160 ;
        RECT 4.000 2254.560 606.000 2334.760 ;
        RECT 4.400 2253.160 606.000 2254.560 ;
        RECT 4.000 2172.960 606.000 2253.160 ;
        RECT 4.400 2171.560 606.000 2172.960 ;
        RECT 4.000 2091.360 606.000 2171.560 ;
        RECT 4.400 2089.960 606.000 2091.360 ;
        RECT 4.000 2009.760 606.000 2089.960 ;
        RECT 4.400 2008.360 606.000 2009.760 ;
        RECT 4.000 1928.160 606.000 2008.360 ;
        RECT 4.400 1926.760 606.000 1928.160 ;
        RECT 4.000 1846.560 606.000 1926.760 ;
        RECT 4.400 1845.160 606.000 1846.560 ;
        RECT 4.000 1764.960 606.000 1845.160 ;
        RECT 4.400 1763.560 606.000 1764.960 ;
        RECT 4.000 1683.360 606.000 1763.560 ;
        RECT 4.400 1681.960 606.000 1683.360 ;
        RECT 4.000 1601.760 606.000 1681.960 ;
        RECT 4.400 1600.360 606.000 1601.760 ;
        RECT 4.000 1520.160 606.000 1600.360 ;
        RECT 4.400 1518.760 606.000 1520.160 ;
        RECT 4.000 1438.560 606.000 1518.760 ;
        RECT 4.400 1437.160 606.000 1438.560 ;
        RECT 4.000 1356.960 606.000 1437.160 ;
        RECT 4.400 1355.560 606.000 1356.960 ;
        RECT 4.000 1275.360 606.000 1355.560 ;
        RECT 4.400 1273.960 606.000 1275.360 ;
        RECT 4.000 1193.760 606.000 1273.960 ;
        RECT 4.400 1192.360 606.000 1193.760 ;
        RECT 4.000 1112.160 606.000 1192.360 ;
        RECT 4.400 1110.760 606.000 1112.160 ;
        RECT 4.000 1030.560 606.000 1110.760 ;
        RECT 4.400 1029.160 606.000 1030.560 ;
        RECT 4.000 948.960 606.000 1029.160 ;
        RECT 4.400 947.560 606.000 948.960 ;
        RECT 4.000 867.360 606.000 947.560 ;
        RECT 4.400 865.960 606.000 867.360 ;
        RECT 4.000 785.760 606.000 865.960 ;
        RECT 4.400 784.360 606.000 785.760 ;
        RECT 4.000 704.160 606.000 784.360 ;
        RECT 4.400 702.760 606.000 704.160 ;
        RECT 4.000 622.560 606.000 702.760 ;
        RECT 4.400 621.160 606.000 622.560 ;
        RECT 4.000 540.960 606.000 621.160 ;
        RECT 4.400 539.560 606.000 540.960 ;
        RECT 4.000 459.360 606.000 539.560 ;
        RECT 4.400 457.960 606.000 459.360 ;
        RECT 4.000 377.760 606.000 457.960 ;
        RECT 4.400 376.360 606.000 377.760 ;
        RECT 4.000 296.160 606.000 376.360 ;
        RECT 4.400 294.760 606.000 296.160 ;
        RECT 4.000 214.560 606.000 294.760 ;
        RECT 4.400 213.160 606.000 214.560 ;
        RECT 4.000 132.960 606.000 213.160 ;
        RECT 4.400 131.560 606.000 132.960 ;
        RECT 4.000 124.800 606.000 131.560 ;
        RECT 4.000 123.400 605.600 124.800 ;
        RECT 4.000 78.560 606.000 123.400 ;
        RECT 4.000 77.160 605.600 78.560 ;
        RECT 4.000 51.360 606.000 77.160 ;
        RECT 4.400 49.960 606.000 51.360 ;
        RECT 4.000 32.320 606.000 49.960 ;
        RECT 4.000 30.920 605.600 32.320 ;
        RECT 4.000 9.015 606.000 30.920 ;
      LAYER met4 ;
        RECT 112.535 11.735 142.240 809.705 ;
        RECT 146.240 11.735 183.040 809.705 ;
        RECT 187.040 11.735 223.840 809.705 ;
        RECT 227.840 11.735 264.640 809.705 ;
        RECT 268.640 11.735 305.440 809.705 ;
        RECT 309.440 11.735 346.240 809.705 ;
        RECT 350.240 11.735 387.040 809.705 ;
        RECT 391.040 11.735 421.985 809.705 ;
  END
END caravel_ips
END LIBRARY

